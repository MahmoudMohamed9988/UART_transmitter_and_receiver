package pkg_receiver;

import uvm_pkg::*;

`include "uvm_macros.svh"
`include "UART_receiver_seq_item.sv"
`include "UART_receiver_sqr.sv"
`include "UART_receiver_agt_config.sv"
`include "UART_receiver_env_config.sv"
`include "UART_receiver_seq.sv"
`include "UART_receiver_vseq.sv"
`include "UART_receiver_drv.sv"
`include "UART_receiver_mon.sv"
`include "UART_receiver_agt.sv"
`include "UART_receiver_evaluator.sv"
`include "UART_receiver_predictor.sv"
`include "UART_receiver_scb.sv"
`include "UART_receiver_cov.sv"
`include "UART_receiver_env.sv"
`include "UART_receiver_test.sv"


endpackage

